//const counter
localparam ZERO8									= 8'd0;
localparam ONE8									= 8'd1;
localparam RAND8									= 8'h0F;
localparam COUNT_MAX4							= 4'd7;