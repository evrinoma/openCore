module MY_NOT(output OUT, input IN);
assign OUT = ~IN;
endmodule
